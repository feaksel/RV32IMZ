// Generated from: factorial.bin
// Total words: 60

imem[  0] = 32'hfd010113;  // addr 0x0000
imem[  1] = 32'h02112623;  // addr 0x0004
imem[  2] = 32'h02812423;  // addr 0x0008
imem[  3] = 32'h03010413;  // addr 0x000c
imem[  4] = 32'hfca42e23;  // addr 0x0010
imem[  5] = 32'hfcb42c23;  // addr 0x0014
imem[  6] = 32'hfe042623;  // addr 0x0018
imem[  7] = 32'hfe042423;  // addr 0x001c
imem[  8] = 32'h0200006f;  // addr 0x0020
imem[  9] = 32'hfec42703;  // addr 0x0024
imem[ 10] = 32'hfdc42783;  // addr 0x0028
imem[ 11] = 32'h00f707b3;  // addr 0x002c
imem[ 12] = 32'hfef42623;  // addr 0x0030
imem[ 13] = 32'hfe842783;  // addr 0x0034
imem[ 14] = 32'h00178793;  // addr 0x0038
imem[ 15] = 32'hfef42423;  // addr 0x003c
imem[ 16] = 32'hfe842783;  // addr 0x0040
imem[ 17] = 32'hfd842703;  // addr 0x0044
imem[ 18] = 32'hfce7cee3;  // addr 0x0048
imem[ 19] = 32'hfec42783;  // addr 0x004c
imem[ 20] = 32'h00078513;  // addr 0x0050
imem[ 21] = 32'h02c12083;  // addr 0x0054
imem[ 22] = 32'h02812403;  // addr 0x0058
imem[ 23] = 32'h03010113;  // addr 0x005c
imem[ 24] = 32'h00008067;  // addr 0x0060
imem[ 25] = 32'hfd010113;  // addr 0x0064
imem[ 26] = 32'h02112623;  // addr 0x0068
imem[ 27] = 32'h02812423;  // addr 0x006c
imem[ 28] = 32'h03010413;  // addr 0x0070
imem[ 29] = 32'hfca42e23;  // addr 0x0074
imem[ 30] = 32'h00100793;  // addr 0x0078
imem[ 31] = 32'hfef42623;  // addr 0x007c
imem[ 32] = 32'hfdc42783;  // addr 0x0080
imem[ 33] = 32'hfef42423;  // addr 0x0084
imem[ 34] = 32'h02c0006f;  // addr 0x0088
imem[ 35] = 32'hfec42783;  // addr 0x008c
imem[ 36] = 32'hfe842703;  // addr 0x0090
imem[ 37] = 32'h00070593;  // addr 0x0094
imem[ 38] = 32'h00078513;  // addr 0x0098
imem[ 39] = 32'hf65ff0ef;  // addr 0x009c
imem[ 40] = 32'h00050793;  // addr 0x00a0
imem[ 41] = 32'hfef42623;  // addr 0x00a4
imem[ 42] = 32'hfe842783;  // addr 0x00a8
imem[ 43] = 32'hfff78793;  // addr 0x00ac
imem[ 44] = 32'hfef42423;  // addr 0x00b0
imem[ 45] = 32'hfe842703;  // addr 0x00b4
imem[ 46] = 32'h00100793;  // addr 0x00b8
imem[ 47] = 32'hfce7c8e3;  // addr 0x00bc
imem[ 48] = 32'hfec42783;  // addr 0x00c0
imem[ 49] = 32'h00078513;  // addr 0x00c4
imem[ 50] = 32'h02c12083;  // addr 0x00c8
imem[ 51] = 32'h02812403;  // addr 0x00cc
imem[ 52] = 32'h03010113;  // addr 0x00d0
imem[ 53] = 32'h00008067;  // addr 0x00d4
imem[ 54] = 32'h00500513;  // addr 0x00d8
imem[ 55] = 32'hf89ff0ef;  // addr 0x00dc
imem[ 56] = 32'h00050793;  // addr 0x00e0
imem[ 57] = 32'h00078513;  // addr 0x00e4
imem[ 58] = 32'h00000013;  // addr 0x00e8
imem[ 59] = 32'hffdff06f;  // addr 0x00ec