// Generated from: factorial_simple.bin
// Total words: 15

imem[  0] = 32'h00100513;  // addr 0x0000
imem[  1] = 32'h00500593;  // addr 0x0004
imem[  2] = 32'h00100293;  // addr 0x0008
imem[  3] = 32'h02b2d463;  // addr 0x000c
imem[  4] = 32'h00050313;  // addr 0x0010
imem[  5] = 32'h00000513;  // addr 0x0014
imem[  6] = 32'h00058393;  // addr 0x0018
imem[  7] = 32'h00038863;  // addr 0x001c
imem[  8] = 32'h00650533;  // addr 0x0020
imem[  9] = 32'hfff38393;  // addr 0x0024
imem[ 10] = 32'hff5ff06f;  // addr 0x0028
imem[ 11] = 32'hfff58593;  // addr 0x002c
imem[ 12] = 32'hfd9ff06f;  // addr 0x0030
imem[ 13] = 32'h0000006f;  // addr 0x0034
imem[ 14] = 32'h00000013;  // addr 0x0038