/**
 * @file tb_c_factorial.v
 * @brief Testbench for factorial program compiled from C
 *
 * Tests the Phase 3 milestone using real compiled C code instead of
 * hand-written assembly. This validates the core against GCC-generated
 * RV32I instructions.
 *
 * Program: factorial(5) = 120
 * Tests: Function calls, loops, branches, stack operations
 *
 * @author RISC-V Core Project
 * @date 2025-12-08
 */

`timescale 1ns / 1ps

module tb_c_factorial;

    reg clk, rst_n;
    initial begin
        clk = 0;
        forever #10 clk = ~clk;
    end

    wire [31:0] iwb_adr_o, iwb_dat_i, dwb_adr_o, dwb_dat_o, dwb_dat_i;
    wire iwb_cyc_o, iwb_stb_o, iwb_ack_i;
    wire dwb_we_o, dwb_cyc_o, dwb_stb_o, dwb_ack_i, dwb_err_i;
    wire [3:0] dwb_sel_o;
    wire [31:0] interrupts;
    assign interrupts = 32'h0;

    // Core with reset vector at address 0
    custom_riscv_core #(
        .RESET_VECTOR(32'h00000000)  // _start at address 0
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        .iwb_adr_o(iwb_adr_o),
        .iwb_dat_i(iwb_dat_i),
        .iwb_cyc_o(iwb_cyc_o),
        .iwb_stb_o(iwb_stb_o),
        .iwb_ack_i(iwb_ack_i),
        .dwb_adr_o(dwb_adr_o),
        .dwb_dat_o(dwb_dat_o),
        .dwb_dat_i(dwb_dat_i),
        .dwb_we_o(dwb_we_o),
        .dwb_sel_o(dwb_sel_o),
        .dwb_cyc_o(dwb_cyc_o),
        .dwb_stb_o(dwb_stb_o),
        .dwb_ack_i(dwb_ack_i),
        .dwb_err_i(dwb_err_i),
        .interrupts(interrupts)
    );

    reg [31:0] imem [0:255];
    reg        imem_ack;
    reg [31:0] dmem [0:255];
    reg        dmem_ack;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            imem_ack <= 1'b0;
        end else begin
            imem_ack <= (iwb_cyc_o && iwb_stb_o && !imem_ack) ? 1'b1 : 1'b0;
        end
    end

    assign iwb_dat_i = (iwb_adr_o[31:2] < 256) ? imem[iwb_adr_o[31:2]] : 32'h00000013;
    assign iwb_ack_i = imem_ack;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            dmem_ack <= 1'b0;
        end else begin
            if (dwb_cyc_o && dwb_stb_o && !dmem_ack) begin
                dmem_ack <= 1'b1;
                if (dwb_we_o && dwb_adr_o[31:2] < 256) begin
                    if (dwb_sel_o[0]) dmem[dwb_adr_o[31:2]][7:0]   <= dwb_dat_o[7:0];
                    if (dwb_sel_o[1]) dmem[dwb_adr_o[31:2]][15:8]  <= dwb_dat_o[15:8];
                    if (dwb_sel_o[2]) dmem[dwb_adr_o[31:2]][23:16] <= dwb_dat_o[23:16];
                    if (dwb_sel_o[3]) dmem[dwb_adr_o[31:2]][31:24] <= dwb_dat_o[31:24];
                end
            end else begin
                dmem_ack <= 1'b0;
            end
        end
    end

    assign dwb_dat_i = (dwb_adr_o[31:2] < 256) ? dmem[dwb_adr_o[31:2]] : 32'h00000000;
    assign dwb_ack_i = dmem_ack;
    assign dwb_err_i = 1'b0;

    integer init_i;

    initial begin
        /**
         * Load compiled C program
         * Generated by: riscv32-unknown-elf-gcc -march=rv32i -O0
         * Source: factorial.c
         */

        // Load program from compiled binary
`include "../../programs/factorial_simple_imem.vh"

        // Fill rest with NOPs
        for (init_i = 15; init_i < 256; init_i = init_i + 1) begin
            imem[init_i] = 32'h00000013;
        end

        // Initialize data memory to zeros
        for (init_i = 0; init_i < 256; init_i = init_i + 1) begin
            dmem[init_i] = 32'h00000000;
        end
    end

    initial begin
        $dumpfile("build/c_factorial.vcd");
        $dumpvars(0, tb_c_factorial);

        rst_n = 0;
        #50;
        rst_n = 1;

        $display("");
        $display("========================================================================");
        $display("PHASE 3 MILESTONE: Factorial from Compiled C Code");
        $display("========================================================================");
        $display("");
        $display("Program: Compiled from C using GCC for RV32I");
        $display("Tests: Function calls (JAL/JALR), loops, branches, stack operations");
        $display("Expected: factorial(5) = 120 in register a0 (x10)");
        $display("");
        $display("Running program...");
        $display("");

        // Run for enough time to complete factorial calculation
        // C code with function calls needs more cycles than hand-written asm
        #100000;

        $display("");
        $display("========================================================================");
        $display("Results");
        $display("========================================================================");
        $display("");
        $display("Return value (a0/x10): %0d (expected: 120)", dut.regfile_inst.registers[10]);
        $display("Stack pointer (sp/x2): 0x%h", dut.regfile_inst.registers[2]);
        $display("Return addr (ra/x1): 0x%h", dut.regfile_inst.registers[1]);
        $display("");

        if (dut.regfile_inst.registers[10] == 32'd120) begin
            $display("*** PHASE 3 MILESTONE PASSED! ***");
            $display("");
            $display("Your core successfully executed:");
            $display("  - GCC-generated RV32I code");
            $display("  - Function calls (JAL/JALR)");
            $display("  - Nested loops");
            $display("  - Conditional branches");
            $display("  - Stack operations (SW/LW with SP)");
            $display("");
            $display("Factorial(5) = %0d (CORRECT!)", dut.regfile_inst.registers[10]);
        end else begin
            $display("*** MILESTONE INCOMPLETE ***");
            $display("");
            $display("Expected factorial(5) = 120");
            $display("Got: %0d", dut.regfile_inst.registers[10]);
            $display("");
            $display("Debug information:");
            $display("  Current PC: 0x%h", dut.pc);
            $display("  a0 (x10) = %0d", dut.regfile_inst.registers[10]);
            $display("  sp (x2)  = 0x%h", dut.regfile_inst.registers[2]);
            $display("  ra (x1)  = 0x%h", dut.regfile_inst.registers[1]);
        end

        $display("========================================================================");
        $display("");

        $finish;
    end

    initial begin
        #200000;
        $display("");
        $display("ERROR: Timeout! Program did not complete in time.");
        $display("This may indicate an infinite loop or stall.");
        $display("Last PC: 0x%h", dut.pc);
        $display("");
        $finish;
    end

endmodule
