# SKY130 LEF (Library Exchange Format) File
# Physical information for standard cells

VERSION 5.8 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

# Technology layers
LAYER met1
  TYPE ROUTING ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  DIRECTION HORIZONTAL ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 0.0361e-3 ;
END met1

LAYER met2  
  TYPE ROUTING ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  DIRECTION VERTICAL ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 0.0200e-3 ;
END met2

LAYER via
  TYPE CUT ;
  SPACING 0.17 ;
  RESISTANCE 4.5 ;
END via

# Standard cell site
SITE unithd
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

# Standard cell definitions
MACRO sky130_fd_sc_hd__inv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.92 BY 2.72 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
      RECT 0.145 0.995 0.315 1.325 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
      RECT 0.605 0.995 0.775 1.325 ;
    END
  END Y
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
      RECT 0 2.480 0.92 2.720 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
      RECT 0 0 0.92 0.240 ;
    END
  END VGND
END sky130_fd_sc_hd__inv_1

MACRO sky130_fd_sc_hd__buf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.84 BY 2.72 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
      RECT 0.145 0.995 0.315 1.325 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
      RECT 1.525 0.995 1.695 1.325 ;
    END
  END X
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
      RECT 0 2.480 1.84 2.720 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
      RECT 0 0 1.84 0.240 ;
    END
  END VGND
END sky130_fd_sc_hd__buf_1

MACRO sky130_fd_sc_hd__dfxtp_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 5.52 BY 2.72 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
      RECT 1.035 0.995 1.205 1.325 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
      RECT 0.145 0.995 0.315 1.325 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
      RECT 5.205 0.995 5.375 1.325 ;
    END
  END Q
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
      RECT 0 2.480 5.52 2.720 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
      RECT 0 0 5.52 0.240 ;
    END
  END VGND
END sky130_fd_sc_hd__dfxtp_1

END LIBRARY