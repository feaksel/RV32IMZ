/**
 * @file tb_c_memory.v
 * @brief Testbench for memory access program compiled from C
 *
 * Tests the Phase 4 milestone using real compiled C code that exercises
 * all load/store operations: LW/SW, LH/SH, LB/SB
 *
 * Program: Memory test with word, halfword, and byte access
 * Tests: Load/store operations, Wishbone bus interface, memory arbiter
 * Expected: sum = 15 + 171 + 10 = 196 in register a0 (x10)
 *
 * @author RISC-V Core Project
 * @date 2025-12-08
 */

`timescale 1ns / 1ps

module tb_c_memory;

    reg clk, rst_n;
    initial begin
        clk = 0;
        forever #10 clk = ~clk;
    end

    wire [31:0] iwb_adr_o, iwb_dat_i, dwb_adr_o, dwb_dat_o, dwb_dat_i;
    wire iwb_cyc_o, iwb_stb_o, iwb_ack_i;
    wire dwb_we_o, dwb_cyc_o, dwb_stb_o, dwb_ack_i, dwb_err_i;
    wire [3:0] dwb_sel_o;
    wire [31:0] interrupts;
    assign interrupts = 32'h0;

    // Core with reset vector at address 0
    custom_riscv_core #(
        .RESET_VECTOR(32'h00000000)
    ) dut (
        .clk(clk),
        .rst_n(rst_n),
        .iwb_adr_o(iwb_adr_o),
        .iwb_dat_i(iwb_dat_i),
        .iwb_cyc_o(iwb_cyc_o),
        .iwb_stb_o(iwb_stb_o),
        .iwb_ack_i(iwb_ack_i),
        .dwb_adr_o(dwb_adr_o),
        .dwb_dat_o(dwb_dat_o),
        .dwb_dat_i(dwb_dat_i),
        .dwb_we_o(dwb_we_o),
        .dwb_sel_o(dwb_sel_o),
        .dwb_cyc_o(dwb_cyc_o),
        .dwb_stb_o(dwb_stb_o),
        .dwb_ack_i(dwb_ack_i),
        .dwb_err_i(dwb_err_i),
        .interrupts(interrupts)
    );

    reg [31:0] imem [0:255];
    reg        imem_ack;
    reg [31:0] dmem [0:255];
    reg        dmem_ack;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            imem_ack <= 1'b0;
        end else begin
            imem_ack <= (iwb_cyc_o && iwb_stb_o && !imem_ack) ? 1'b1 : 1'b0;
        end
    end

    assign iwb_dat_i = (iwb_adr_o[31:2] < 256) ? imem[iwb_adr_o[31:2]] : 32'h00000013;
    assign iwb_ack_i = imem_ack;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            dmem_ack <= 1'b0;
        end else begin
            if (dwb_cyc_o && dwb_stb_o && !dmem_ack) begin
                dmem_ack <= 1'b1;
                if (dwb_we_o && dwb_adr_o[31:2] < 256) begin
                    if (dwb_sel_o[0]) dmem[dwb_adr_o[31:2]][7:0]   <= dwb_dat_o[7:0];
                    if (dwb_sel_o[1]) dmem[dwb_adr_o[31:2]][15:8]  <= dwb_dat_o[15:8];
                    if (dwb_sel_o[2]) dmem[dwb_adr_o[31:2]][23:16] <= dwb_dat_o[23:16];
                    if (dwb_sel_o[3]) dmem[dwb_adr_o[31:2]][31:24] <= dwb_dat_o[31:24];
                end
            end else begin
                dmem_ack <= 1'b0;
            end
        end
    end

    assign dwb_dat_i = (dwb_adr_o[31:2] < 256) ? dmem[dwb_adr_o[31:2]] : 32'h00000000;
    assign dwb_ack_i = dmem_ack;
    assign dwb_err_i = 1'b0;

    integer init_i;

    initial begin
        /**
         * Load compiled C program
         * Generated by: riscv32-unknown-elf-gcc -march=rv32i
         * Source: memory_test.c
         */

        // Load program from compiled binary
`include "../../programs/memory_test_imem.vh"

        // Fill rest with NOPs
        for (init_i = 34; init_i < 256; init_i = init_i + 1) begin
            imem[init_i] = 32'h00000013;
        end

        // Initialize data memory to zeros
        for (init_i = 0; init_i < 256; init_i = init_i + 1) begin
            dmem[init_i] = 32'h00000000;
        end
    end

    initial begin
        $dumpfile("build/c_memory.vcd");
        $dumpvars(0, tb_c_memory);

        rst_n = 0;
        #50;
        rst_n = 1;

        $display("");
        $display("========================================================================");
        $display("PHASE 4 MILESTONE: Memory Access from Compiled C Code");
        $display("========================================================================");
        $display("");
        $display("Program: Compiled from C using GCC for RV32I");
        $display("Tests: Word/Halfword/Byte Load/Store, Wishbone bus interface");
        $display("");
        $display("Operations:");
        $display("  1. Store words: 1, 2, 3, 4, 5 (SW)");
        $display("  2. Load words and sum (LW)");
        $display("  3. Store and load halfword: 0xAB = 171 (SH/LH)");
        $display("  4. Store and load byte: 10 (SB/LB)");
        $display("");
        $display("Expected result: 1+2+3+4+5+171+10 = 196 in a0");
        $display("");
        $display("Running program...");
        $display("");

        // Run for enough time to complete memory operations
        #10000;

        $display("");
        $display("========================================================================");
        $display("Results");
        $display("========================================================================");
        $display("");
        $display("Result (a0/x10): %0d (expected: 196)", dut.regfile_inst.registers[10]);
        $display("");

        // Check memory contents
        $display("Data Memory Contents:");
        $display("  dmem[0x40] (word 64, addr 0x100): 0x%h (expected: 0x00000001)", dmem[64]);
        $display("  dmem[0x41] (word 65, addr 0x104): 0x%h (expected: 0x00000002)", dmem[65]);
        $display("  dmem[0x42] (word 66, addr 0x108): 0x%h (expected: 0x00000003)", dmem[66]);
        $display("  dmem[0x43] (word 67, addr 0x10C): 0x%h (expected: 0x00000004)", dmem[67]);
        $display("  dmem[0x44] (word 68, addr 0x110): 0x%h (expected: 0x00000005)", dmem[68]);
        $display("  dmem[0x48] (word 72, addr 0x120): 0x%h (expected: 0x000000AB halfword)", dmem[72]);
        $display("  dmem[0x4C] (word 76, addr 0x130): 0x%h (expected: 0x0000000A byte)", dmem[76]);
        $display("");

        if (dut.regfile_inst.registers[10] == 32'd196 &&
            dmem[64] == 32'd1 &&
            dmem[65] == 32'd2 &&
            dmem[66] == 32'd3 &&
            dmem[67] == 32'd4 &&
            dmem[68] == 32'd5 &&
            (dmem[72] & 32'h0000FFFF) == 32'h000000AB &&
            (dmem[76] & 32'h000000FF) == 32'h0000000A) begin
            $display("*** PHASE 4 MILESTONE PASSED! ***");
            $display("");
            $display("Your core successfully executed:");
            $display("  - Word load/store (LW/SW)");
            $display("  - Halfword load/store (LH/SH)");
            $display("  - Byte load/store (LB/SB)");
            $display("  - Wishbone bus transactions");
            $display("  - Byte-select write operations");
            $display("");
            $display("Memory result = %0d (CORRECT!)", dut.regfile_inst.registers[10]);
        end else begin
            $display("*** MILESTONE INCOMPLETE ***");
            $display("");
            $display("Expected result = 196");
            $display("Got: %0d", dut.regfile_inst.registers[10]);
            $display("");
            $display("Debug information:");
            $display("  Current PC: 0x%h", dut.pc);
            $display("  a0 (x10) = %0d", dut.regfile_inst.registers[10]);
            $display("  a1 (x11) = 0x%h (base addr)", dut.regfile_inst.registers[11]);
        end

        $display("========================================================================");
        $display("");

        $finish;
    end

    initial begin
        #50000;
        $display("");
        $display("ERROR: Timeout! Program did not complete in time.");
        $display("Last PC: 0x%h", dut.pc);
        $display("");
        $finish;
    end

endmodule
