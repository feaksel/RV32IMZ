module test_syntax;\n    // Just instantiate the core to test syntax\n    \n    wire clk = 1'b0;\n    wire rst_n = 1'b1;\n    \n    custom_riscv_core core (\n        .clk(clk),\n        .rst_n(rst_n),\n        .iwb_adr_o(),\n        .iwb_dat_i(32'h0),\n        .iwb_cyc_o(),\n        .iwb_stb_o(),\n        .iwb_ack_i(1'b0),\n        .iwb_err_i(1'b0),\n        .dwb_adr_o(),\n        .dwb_dat_o(),\n        .dwb_dat_i(32'h0),\n        .dwb_we_o(),\n        .dwb_sel_o(),\n        .dwb_cyc_o(),\n        .dwb_stb_o(),\n        .dwb_ack_i(1'b0),\n        .dwb_err_i(1'b0),\n        .interrupts(32'h0)\n    );\n    \nendmodule\n