// Generated from: memory_test.bin
// Total words: 34

imem[  0] = 32'h10000593;  // addr 0x0000
imem[  1] = 32'h00100293;  // addr 0x0004
imem[  2] = 32'h0055a023;  // addr 0x0008
imem[  3] = 32'h00200293;  // addr 0x000c
imem[  4] = 32'h0055a223;  // addr 0x0010
imem[  5] = 32'h00300293;  // addr 0x0014
imem[  6] = 32'h0055a423;  // addr 0x0018
imem[  7] = 32'h00400293;  // addr 0x001c
imem[  8] = 32'h0055a623;  // addr 0x0020
imem[  9] = 32'h00500293;  // addr 0x0024
imem[ 10] = 32'h0055a823;  // addr 0x0028
imem[ 11] = 32'h00000513;  // addr 0x002c
imem[ 12] = 32'h0005a303;  // addr 0x0030
imem[ 13] = 32'h00650533;  // addr 0x0034
imem[ 14] = 32'h0045a303;  // addr 0x0038
imem[ 15] = 32'h00650533;  // addr 0x003c
imem[ 16] = 32'h0085a303;  // addr 0x0040
imem[ 17] = 32'h00650533;  // addr 0x0044
imem[ 18] = 32'h00c5a303;  // addr 0x0048
imem[ 19] = 32'h00650533;  // addr 0x004c
imem[ 20] = 32'h0105a303;  // addr 0x0050
imem[ 21] = 32'h00650533;  // addr 0x0054
imem[ 22] = 32'h12000613;  // addr 0x0058
imem[ 23] = 32'h0ab00293;  // addr 0x005c
imem[ 24] = 32'h00561023;  // addr 0x0060
imem[ 25] = 32'h00061303;  // addr 0x0064
imem[ 26] = 32'h00650533;  // addr 0x0068
imem[ 27] = 32'h13000693;  // addr 0x006c
imem[ 28] = 32'h00a00293;  // addr 0x0070
imem[ 29] = 32'h00568023;  // addr 0x0074
imem[ 30] = 32'h00068303;  // addr 0x0078
imem[ 31] = 32'h00650533;  // addr 0x007c
imem[ 32] = 32'h0000006f;  // addr 0x0080
imem[ 33] = 32'h00000013;  // addr 0x0084