# SKY130 Technology LEF File
# Physical technology information

VERSION 5.8 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

# Process technology layers
LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER diff
  TYPE MASTERSLICE ;
END diff

LAYER tap
  TYPE MASTERSLICE ;
END tap

LAYER poly
  TYPE MASTERSLICE ;
END poly

LAYER licon1
  TYPE CUT ;
  SPACING 0.17 ;
END licon1

LAYER li1
  TYPE ROUTING ;
  PITCH 0.48 ;
  WIDTH 0.17 ;
  SPACING 0.17 ;
  RESISTANCE RPERSQ 12.2 ;
END li1

LAYER mcon
  TYPE CUT ;
  SPACING 0.19 ;
END mcon

LAYER met1
  TYPE ROUTING ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  DIRECTION HORIZONTAL ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 0.0361e-3 ;
  EDGECAPACITANCE 0.0281e-6 ;
END met1

LAYER via
  TYPE CUT ;
  SPACING 0.17 ;
  RESISTANCE 4.5 ;
END via

LAYER met2
  TYPE ROUTING ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
  SPACING 0.14 ;
  DIRECTION VERTICAL ;
  RESISTANCE RPERSQ 0.125 ;
  CAPACITANCE CPERSQDIST 0.0200e-3 ;
  EDGECAPACITANCE 0.0281e-6 ;
END met2

LAYER via2
  TYPE CUT ;
  SPACING 0.20 ;
  RESISTANCE 4.5 ;
END via2

LAYER met3
  TYPE ROUTING ;
  PITCH 0.68 ;
  WIDTH 0.30 ;
  SPACING 0.30 ;
  DIRECTION HORIZONTAL ;
  RESISTANCE RPERSQ 0.047 ;
  CAPACITANCE CPERSQDIST 0.0136e-3 ;
  EDGECAPACITANCE 0.0281e-6 ;
END met3

LAYER via3
  TYPE CUT ;
  SPACING 0.20 ;
  RESISTANCE 4.5 ;
END via3

LAYER met4
  TYPE ROUTING ;
  PITCH 0.92 ;
  WIDTH 0.30 ;
  SPACING 0.30 ;
  DIRECTION VERTICAL ;
  RESISTANCE RPERSQ 0.047 ;
  CAPACITANCE CPERSQDIST 0.0103e-3 ;
  EDGECAPACITANCE 0.0281e-6 ;
END met4

LAYER via4
  TYPE CUT ;
  SPACING 0.20 ;
  RESISTANCE 4.5 ;
END via4

LAYER met5
  TYPE ROUTING ;
  PITCH 3.44 ;
  WIDTH 1.60 ;
  SPACING 1.60 ;
  DIRECTION HORIZONTAL ;
  RESISTANCE RPERSQ 0.029 ;
  CAPACITANCE CPERSQDIST 0.0074e-3 ;
  EDGECAPACITANCE 0.0281e-6 ;
END met5

# Standard cell site
SITE unithd
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

END LIBRARY